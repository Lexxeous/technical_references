--VHDL Coding Reference